library verilog;
use verilog.vl_types.all;
entity computer_vlg_vec_tst is
end computer_vlg_vec_tst;
