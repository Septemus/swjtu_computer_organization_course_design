library verilog;
use verilog.vl_types.all;
entity reg_function_vlg_vec_tst is
end reg_function_vlg_vec_tst;
